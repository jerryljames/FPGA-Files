`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:33:52 12/12/2014 
// Design Name: 
// Module Name:    Synchronous_Up_Down_Counter_74HC193 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 5.	Design a 4-Bit synchronous up/down counter (dual clock with clear).  Refer datasheet of 74HC193 for the detailed functional description
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Synchronous_Up_Down_Counter_74HC193(CPU,CPD,MR,Q,D,PL_BAR);
input CPU,CPD,MR,PL_BAR;
input [3:0]D;
output [3:0]Q;
always @(CPD)



endmodule
